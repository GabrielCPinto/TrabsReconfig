library ieee;
use ieee.std_logic_1164.all;

ENTITY control_unity IS
	PORT(
		nrst			: IN STD_LOGIC;		
		clk				: IN STD_LOGIC;		
		instr			: IN STD_LOGIC_VECTOR(13 DOWNTO 0);
		alu_z			: IN STD_LOGIC;

		op_sel 			: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		bit_sel			: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		wr_z_en			: OUT STD_LOGIC;
		wr_dc_en		: OUT STD_LOGIC;
		wr_c_en			: OUT STD_LOGIC;
		wr_w_reg_en		: OUT STD_LOGIC;
		wr_en			: OUT STD_LOGIC;
		rd_en			: OUT STD_LOGIC;
		load_pc			: OUT STD_LOGIC;
		inc_pc			: OUT STD_LOGIC;
		stack_push		: OUT STD_LOGIC;
		stack_pop		: OUT STD_LOGIC;
		lit_sel			: OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE arch1 OF control_unity IS
	TYPE state_type IS (rst, fetch_only, fet_dec_ex);
	SIGNAL pres_state 	: state_type;	
	SIGNAL next_state 	: state_type;

	---------BYTE-ORIENTED FILE REGISTER OPERATIONS--------------------------------

	CONSTANT ADDWF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000111";
	CONSTANT ANDWF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000101";
	CONSTANT CLRF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000001";
	CONSTANT CLRW		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000001";
	CONSTANT COMF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "001001";
	CONSTANT DECF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000011";
	CONSTANT DECFSZ		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "001011";
	CONSTANT INCF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "001010";
	CONSTANT INCFSZ		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "001111";
	CONSTANT IORWF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000100";
	CONSTANT MOVF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "001000";
	CONSTANT MOVWF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000000";
	CONSTANT NOP		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000000";
	CONSTANT RLF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "001101";
	CONSTANT RRF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "001100";
	CONSTANT SUBWF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000010";
	CONSTANT SWAPF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "001110";
	CONSTANT XORWF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000110";

	------BIT-ORIENTED FILE REGISTER OPERATIONS-------------------------

	CONSTANT BCF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "0100";
	CONSTANT BSF		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "0101";
	CONSTANT BTFSC		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "0110";
	CONSTANT BTFSS		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "0111";

	-------LITERAL AND CONTROL OPERATIONS----------------------------
	CONSTANT ADDLW		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "11111";
	CONSTANT ANDLW		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "111001";
	CONSTANT CALL		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "100";
	CONSTANT CLRWDT		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000000";
	CONSTANT GOTO		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "101";
	CONSTANT IORLW		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "111000";
	CONSTANT MOVLW		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "1100";
	CONSTANT RETFIE		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000000";
	CONSTANT RETLW		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "1101";
	CONSTANT RET_URN	: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000000";
	CONSTANT SLEEP		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "000000";
	CONSTANT SUBLW		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "11110x";
	CONSTANT XORLW		: STD_LOGIC_VECTOR(7 DOWNTO 0) := "111010";

BEGIN

	inc_pc <= '1';
	load_pc
	stack_push
	stack_pop
	bit_sel[2..0] <= "----"
	
	wr_z_en
	wr_dc_en
	wr_c_en
	rd_en
	lit_sel

	case instr is 
	when instr(5 downto 0) = ADDWF =>

	op_sel[3..0] <= codigo de adicionar na ULA

	IF(instruction(6) = '0') THEN 
		wr_w_reg_en <= '1'

	ELSE 
	wr_en <= 1;

--tudo que for registrar F pode assumir q � memoira
--tudo que for regi

END arch1;