LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY RAM_mem IS
PORT (
	nrst : IN STD_LOGIC; --Entrada de reset assíncrono. Quando ativada (nível lógico baixo), todos os bits da memória
--RAM deverão ser zerados. Esta entrada tem preferência sobre todas as outras.
	clk_in : IN STD_LOGIC; --Entrada de clock do sistema. A escrita na memória acontece na borda de subida do clock,
--desde que habilitada.
	wr_en : IN STD_LOGIC; --Entrada de habilitação para escrita na memória. Quando ativada (nível lógico alto), a
--memória será escrita, síncrona com clk_in, com o valor de dbus_in, desde que o endereço correspondente esteja 
--presente em abus_in, conforme especificado no item 3.3. Caso contrário, nenhuma ação será efetuada. 
	rd_en : IN STD_LOGIC; --Entrada de habilitação para leitura. Quando ativada (nível lógico alto), a saída dbus_out
--deverá corresponder ao conteúdo da memória endereçada. Quando desativada ou quando o endereço não corresponder 
--ao especificado no item 3.3, a saída deverá ficar em alta impedância (“ZZZZZZZZ”). 
	abus_in :  IN STD_LOGIC_VECTOR (8 DOWNTO 0); --Entrada de endereçamento. Aponta a célula de memória a ser 
--escrita ou lida, desde que habilitada. As faixas de endereço para cada área de memória estão definidas no item 3.3.
	dbus_in :  IN STD_LOGIC_VECTOR (7 DOWNTO 0); --Entrada de dados para escrita na memória, com habilitação 
--através de wr_en, e endereçamento por abus_in.
	dbus_out :  OUT STD_LOGIC_VECTOR (7 DOWNTO 0) --Barramento de saída de dados, com 8 bits. Habilitação a
--través de rd_en e endereçamento por abus_in. Durante as operações de leitura, comporta-se como saída. 
--Quando não em uso, fica em alta impedância (“ZZZZZZZZ”). A operação de leitura deve ser completamente
--combinacional, ou seja, não depende de transição de clk_in.
);
END ENTITY;

ARCHITECTURE arch1 OF RAM_mem IS
	TYPE memory_type0 IS ARRAY (32 TO 111) OF STD_LOGIC_VECTOR (7 DOWNTO 0); --Array de 80 bytes
	TYPE memory_type1 IS ARRAY (160 TO 239) OF STD_LOGIC_VECTOR (7 DOWNTO 0); --Array de 80 bytes
	TYPE memory_type2 IS ARRAY (288 TO 367) OF STD_LOGIC_VECTOR (7 DOWNTO 0); --Array de 80 bytes
	TYPE small_memory_type IS ARRAY (112 TO 127) OF STD_LOGIC_VECTOR (7 DOWNTO 0);	 --Array 16 bytes
	
	SIGNAL mem0 : memory_type0; --Primeira área de memória
	SIGNAL mem1 : memory_type1; --Segunda área de memória
	SIGNAL mem2 : memory_type2; --Terceira área de memória
	SIGNAL mem_com : small_memory_type; --Quarta área de memória
BEGIN
	PROCESS(nrst, clk_in) 
		BEGIN
		
		IF nrst = '0' THEN  --Limpa toda área da RAM
			FOR i IN 0 TO 79 LOOP --Loop das áreas com 80bytes
				mem0(i) <= (OTHERS => '0'); 
				mem1(i) <= (OTHERS => '0');
				mem2(i) <= (OTHERS => '0');
			END LOOP;
			
			FOR i IN 0 TO 15 LOOP --loop da área com 16bytes
				mem_com(i) <= (OTHERS => '0');
			END LOOP;
			
		ELSIF RISING_EDGE(clk_in) AND wr_en = '1' THEN  --Escrita na memoria de forma sincrona
            
            IF abus_in >= x"20" AND abus_in <= x"6F" THEN --validações da área de memoria selecionada
				mem0(to_integer(unsigned(abus_in))) <= dbus_in; 
            ELSIF abus_in >= x"A0" AND abus_in <= x"EF" THEN --validações da área de memoria selecionada
                mem1(to_integer(unsigned(abus_in))) <= dbus_in; 
            ELSIF abus_in >= x"120" AND abus_in <= x"16F" THEN --validações da área de memoria selecionada
                mem2(to_integer(unsigned(abus_in))) <= dbus_in; 
            ELSIF abus_in >= x"70" AND abus_in <= x"7F" THEN --validações da área de memoria selecionada
                mem_com(to_integer(unsigned(abus_in))) <= dbus_in; 
            END IF;
			
		END IF;
	END PROCESS;

    PROCESS(rd_en)
        BEGIN
        IF rd_en = '0' THEN
            dbus_out <= "ZZZZZZZZ";
        ELSIF rd_en = '1' THEN

            IF abus_in >= x"20" AND abus_in <= x"6F" THEN --validações da área de memoria selecionada
                dbus_out <= mem0(to_integer(unsigned(abus_in))); 
            ELSIF abus_in >= x"A0" AND abus_in <= x"EF" THEN --validações da área de memoria selecionada
                dbus_out <= mem1(to_integer(unsigned(abus_in))); 
            ELSIF abus_in >= x"120" AND abus_in <= x"16F" THEN --validações da área de memoria selecionada
                dbus_out <= mem2(to_integer(unsigned(abus_in))); 
            ELSIF abus_in >= x"70" AND abus_in <= x"7F" THEN --validações da área de memoria selecionada
                dbus_out <= mem_com(to_integer(unsigned(abus_in))); 
            END IF;

        END IF;
    END PROCESS;
END arch1;
